/*
to debugg

in cmd

+access+r+UVM_PHASE_TRACE


*/

