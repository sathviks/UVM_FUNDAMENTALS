/*
to debugg

in cmd

+access+r+UVM_OBJECTION_TRACE


*/


